`define FSM_WIDTH 8 
// `CLP
`define VIVADO_ENV